library ieee;
library work;
use ieee.std_logic_1164;